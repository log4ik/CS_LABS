library verilog;
use verilog.vl_types.all;
entity decoder8_tb is
end decoder8_tb;
