library verilog;
use verilog.vl_types.all;
entity Lohovskyi_lab4 is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        f1              : out    vl_logic;
        f2              : out    vl_logic
    );
end Lohovskyi_lab4;
